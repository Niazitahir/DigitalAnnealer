// DE1_SOC.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module DE1_SOC (
		input  wire        clk_clk,                         //                  clk.clk
		input  wire        hps_0_h2f_mpu_events_eventi,     // hps_0_h2f_mpu_events.eventi
		output wire        hps_0_h2f_mpu_events_evento,     //                     .evento
		output wire [1:0]  hps_0_h2f_mpu_events_standbywfe, //                     .standbywfe
		output wire [1:0]  hps_0_h2f_mpu_events_standbywfi, //                     .standbywfi
		output wire [12:0] memory_mem_a,                    //               memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                     .mem_ba
		output wire        memory_mem_ck,                   //                     .mem_ck
		output wire        memory_mem_ck_n,                 //                     .mem_ck_n
		output wire        memory_mem_cke,                  //                     .mem_cke
		output wire        memory_mem_cs_n,                 //                     .mem_cs_n
		output wire        memory_mem_ras_n,                //                     .mem_ras_n
		output wire        memory_mem_cas_n,                //                     .mem_cas_n
		output wire        memory_mem_we_n,                 //                     .mem_we_n
		output wire        memory_mem_reset_n,              //                     .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                   //                     .mem_dq
		inout  wire        memory_mem_dqs,                  //                     .mem_dqs
		inout  wire        memory_mem_dqs_n,                //                     .mem_dqs_n
		output wire        memory_mem_odt,                  //                     .mem_odt
		output wire        memory_mem_dm,                   //                     .mem_dm
		input  wire        memory_oct_rzqin                 //                     .oct_rzqin
	);

	wire         sys_sdram_pll_0_sdram_clk_clk;                                // sys_sdram_pll_0:sdram_clk_clk -> hps_0:f2h_sdram0_clk
	wire         sys_sdram_pll_0_sys_clk_clk;                                  // sys_sdram_pll_0:sys_clk_clk -> [hps_0:f2h_axi_clk, hps_0:h2f_axi_clk, hps_0:h2f_lw_axi_clk, jtag_uart_0:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, mm_interconnect_1:sys_sdram_pll_0_sys_clk_clk, rst_controller:clk, single_port_ram_0:clk]
	wire         hps_0_h2f_reset_reset;                                        // hps_0:h2f_rst_n -> [rst_controller:reset_in0, sys_sdram_pll_0:ref_reset_reset]
	wire   [1:0] hps_0_h2f_axi_master_awburst;                                 // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                                   // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [7:0] hps_0_h2f_axi_master_wstrb;                                   // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                                  // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                                     // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                                  // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                                   // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                                     // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                                 // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                                  // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                                  // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                                  // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                                  // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [63:0] hps_0_h2f_axi_master_wdata;                                   // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                                 // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                                 // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                                    // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                                  // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                                  // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                                  // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                                   // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                                 // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [63:0] hps_0_h2f_axi_master_rdata;                                   // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                                 // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                                 // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                                  // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                                  // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                                   // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                                   // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                                   // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                                    // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                                     // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                                  // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                                  // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                                 // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                                  // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire   [7:0] mm_interconnect_0_single_port_ram_0_avalon_slave_0_readdata;  // single_port_ram_0:q -> mm_interconnect_0:single_port_ram_0_avalon_slave_0_readdata
	wire   [5:0] mm_interconnect_0_single_port_ram_0_avalon_slave_0_address;   // mm_interconnect_0:single_port_ram_0_avalon_slave_0_address -> single_port_ram_0:addr
	wire         mm_interconnect_0_single_port_ram_0_avalon_slave_0_write;     // mm_interconnect_0:single_port_ram_0_avalon_slave_0_write -> single_port_ram_0:we
	wire   [7:0] mm_interconnect_0_single_port_ram_0_avalon_slave_0_writedata; // mm_interconnect_0:single_port_ram_0_avalon_slave_0_writedata -> single_port_ram_0:data
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                              // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                                // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                                // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                               // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                  // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                               // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                                // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                  // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                              // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                               // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                               // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                               // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                               // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                                // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                              // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                              // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                 // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                               // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                               // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                               // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                                // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                              // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                                // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                              // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                              // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                               // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                               // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                                // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                                // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                                // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                 // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                  // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                               // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                               // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                              // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                               // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [jtag_uart_0:rst_n, mm_interconnect_0:single_port_ram_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_0_reset_reset_bridge_in_reset_reset, single_port_ram_0:reset_n]

	DE1_SOC_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.h2f_mpu_eventi     (hps_0_h2f_mpu_events_eventi),     //    h2f_mpu_events.eventi
		.h2f_mpu_evento     (hps_0_h2f_mpu_events_evento),     //                  .evento
		.h2f_mpu_standbywfe (hps_0_h2f_mpu_events_standbywfe), //                  .standbywfe
		.h2f_mpu_standbywfi (hps_0_h2f_mpu_events_standbywfi), //                  .standbywfi
		.mem_a              (memory_mem_a),                    //            memory.mem_a
		.mem_ba             (memory_mem_ba),                   //                  .mem_ba
		.mem_ck             (memory_mem_ck),                   //                  .mem_ck
		.mem_ck_n           (memory_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke            (memory_mem_cke),                  //                  .mem_cke
		.mem_cs_n           (memory_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n          (memory_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n           (memory_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),              //                  .mem_reset_n
		.mem_dq             (memory_mem_dq),                   //                  .mem_dq
		.mem_dqs            (memory_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt            (memory_mem_odt),                  //                  .mem_odt
		.mem_dm             (memory_mem_dm),                   //                  .mem_dm
		.oct_rzqin          (memory_oct_rzqin),                //                  .oct_rzqin
		.h2f_rst_n          (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.f2h_sdram0_clk     (sys_sdram_pll_0_sdram_clk_clk),   //  f2h_sdram0_clock.clk
		.f2h_sdram0_ARADDR  (),                                //   f2h_sdram0_data.araddr
		.f2h_sdram0_ARLEN   (),                                //                  .arlen
		.f2h_sdram0_ARID    (),                                //                  .arid
		.f2h_sdram0_ARSIZE  (),                                //                  .arsize
		.f2h_sdram0_ARBURST (),                                //                  .arburst
		.f2h_sdram0_ARLOCK  (),                                //                  .arlock
		.f2h_sdram0_ARPROT  (),                                //                  .arprot
		.f2h_sdram0_ARVALID (),                                //                  .arvalid
		.f2h_sdram0_ARCACHE (),                                //                  .arcache
		.f2h_sdram0_AWADDR  (),                                //                  .awaddr
		.f2h_sdram0_AWLEN   (),                                //                  .awlen
		.f2h_sdram0_AWID    (),                                //                  .awid
		.f2h_sdram0_AWSIZE  (),                                //                  .awsize
		.f2h_sdram0_AWBURST (),                                //                  .awburst
		.f2h_sdram0_AWLOCK  (),                                //                  .awlock
		.f2h_sdram0_AWPROT  (),                                //                  .awprot
		.f2h_sdram0_AWVALID (),                                //                  .awvalid
		.f2h_sdram0_AWCACHE (),                                //                  .awcache
		.f2h_sdram0_BRESP   (),                                //                  .bresp
		.f2h_sdram0_BID     (),                                //                  .bid
		.f2h_sdram0_BVALID  (),                                //                  .bvalid
		.f2h_sdram0_BREADY  (),                                //                  .bready
		.f2h_sdram0_ARREADY (),                                //                  .arready
		.f2h_sdram0_AWREADY (),                                //                  .awready
		.f2h_sdram0_RREADY  (),                                //                  .rready
		.f2h_sdram0_RDATA   (),                                //                  .rdata
		.f2h_sdram0_RRESP   (),                                //                  .rresp
		.f2h_sdram0_RLAST   (),                                //                  .rlast
		.f2h_sdram0_RID     (),                                //                  .rid
		.f2h_sdram0_RVALID  (),                                //                  .rvalid
		.f2h_sdram0_WLAST   (),                                //                  .wlast
		.f2h_sdram0_WVALID  (),                                //                  .wvalid
		.f2h_sdram0_WDATA   (),                                //                  .wdata
		.f2h_sdram0_WSTRB   (),                                //                  .wstrb
		.f2h_sdram0_WREADY  (),                                //                  .wready
		.f2h_sdram0_WID     (),                                //                  .wid
		.h2f_axi_clk        (sys_sdram_pll_0_sys_clk_clk),     //     h2f_axi_clock.clk
		.h2f_AWID           (hps_0_h2f_axi_master_awid),       //    h2f_axi_master.awid
		.h2f_AWADDR         (hps_0_h2f_axi_master_awaddr),     //                  .awaddr
		.h2f_AWLEN          (hps_0_h2f_axi_master_awlen),      //                  .awlen
		.h2f_AWSIZE         (hps_0_h2f_axi_master_awsize),     //                  .awsize
		.h2f_AWBURST        (hps_0_h2f_axi_master_awburst),    //                  .awburst
		.h2f_AWLOCK         (hps_0_h2f_axi_master_awlock),     //                  .awlock
		.h2f_AWCACHE        (hps_0_h2f_axi_master_awcache),    //                  .awcache
		.h2f_AWPROT         (hps_0_h2f_axi_master_awprot),     //                  .awprot
		.h2f_AWVALID        (hps_0_h2f_axi_master_awvalid),    //                  .awvalid
		.h2f_AWREADY        (hps_0_h2f_axi_master_awready),    //                  .awready
		.h2f_WID            (hps_0_h2f_axi_master_wid),        //                  .wid
		.h2f_WDATA          (hps_0_h2f_axi_master_wdata),      //                  .wdata
		.h2f_WSTRB          (hps_0_h2f_axi_master_wstrb),      //                  .wstrb
		.h2f_WLAST          (hps_0_h2f_axi_master_wlast),      //                  .wlast
		.h2f_WVALID         (hps_0_h2f_axi_master_wvalid),     //                  .wvalid
		.h2f_WREADY         (hps_0_h2f_axi_master_wready),     //                  .wready
		.h2f_BID            (hps_0_h2f_axi_master_bid),        //                  .bid
		.h2f_BRESP          (hps_0_h2f_axi_master_bresp),      //                  .bresp
		.h2f_BVALID         (hps_0_h2f_axi_master_bvalid),     //                  .bvalid
		.h2f_BREADY         (hps_0_h2f_axi_master_bready),     //                  .bready
		.h2f_ARID           (hps_0_h2f_axi_master_arid),       //                  .arid
		.h2f_ARADDR         (hps_0_h2f_axi_master_araddr),     //                  .araddr
		.h2f_ARLEN          (hps_0_h2f_axi_master_arlen),      //                  .arlen
		.h2f_ARSIZE         (hps_0_h2f_axi_master_arsize),     //                  .arsize
		.h2f_ARBURST        (hps_0_h2f_axi_master_arburst),    //                  .arburst
		.h2f_ARLOCK         (hps_0_h2f_axi_master_arlock),     //                  .arlock
		.h2f_ARCACHE        (hps_0_h2f_axi_master_arcache),    //                  .arcache
		.h2f_ARPROT         (hps_0_h2f_axi_master_arprot),     //                  .arprot
		.h2f_ARVALID        (hps_0_h2f_axi_master_arvalid),    //                  .arvalid
		.h2f_ARREADY        (hps_0_h2f_axi_master_arready),    //                  .arready
		.h2f_RID            (hps_0_h2f_axi_master_rid),        //                  .rid
		.h2f_RDATA          (hps_0_h2f_axi_master_rdata),      //                  .rdata
		.h2f_RRESP          (hps_0_h2f_axi_master_rresp),      //                  .rresp
		.h2f_RLAST          (hps_0_h2f_axi_master_rlast),      //                  .rlast
		.h2f_RVALID         (hps_0_h2f_axi_master_rvalid),     //                  .rvalid
		.h2f_RREADY         (hps_0_h2f_axi_master_rready),     //                  .rready
		.f2h_axi_clk        (sys_sdram_pll_0_sys_clk_clk),     //     f2h_axi_clock.clk
		.f2h_AWID           (),                                //     f2h_axi_slave.awid
		.f2h_AWADDR         (),                                //                  .awaddr
		.f2h_AWLEN          (),                                //                  .awlen
		.f2h_AWSIZE         (),                                //                  .awsize
		.f2h_AWBURST        (),                                //                  .awburst
		.f2h_AWLOCK         (),                                //                  .awlock
		.f2h_AWCACHE        (),                                //                  .awcache
		.f2h_AWPROT         (),                                //                  .awprot
		.f2h_AWVALID        (),                                //                  .awvalid
		.f2h_AWREADY        (),                                //                  .awready
		.f2h_AWUSER         (),                                //                  .awuser
		.f2h_WID            (),                                //                  .wid
		.f2h_WDATA          (),                                //                  .wdata
		.f2h_WSTRB          (),                                //                  .wstrb
		.f2h_WLAST          (),                                //                  .wlast
		.f2h_WVALID         (),                                //                  .wvalid
		.f2h_WREADY         (),                                //                  .wready
		.f2h_BID            (),                                //                  .bid
		.f2h_BRESP          (),                                //                  .bresp
		.f2h_BVALID         (),                                //                  .bvalid
		.f2h_BREADY         (),                                //                  .bready
		.f2h_ARID           (),                                //                  .arid
		.f2h_ARADDR         (),                                //                  .araddr
		.f2h_ARLEN          (),                                //                  .arlen
		.f2h_ARSIZE         (),                                //                  .arsize
		.f2h_ARBURST        (),                                //                  .arburst
		.f2h_ARLOCK         (),                                //                  .arlock
		.f2h_ARCACHE        (),                                //                  .arcache
		.f2h_ARPROT         (),                                //                  .arprot
		.f2h_ARVALID        (),                                //                  .arvalid
		.f2h_ARREADY        (),                                //                  .arready
		.f2h_ARUSER         (),                                //                  .aruser
		.f2h_RID            (),                                //                  .rid
		.f2h_RDATA          (),                                //                  .rdata
		.f2h_RRESP          (),                                //                  .rresp
		.f2h_RLAST          (),                                //                  .rlast
		.f2h_RVALID         (),                                //                  .rvalid
		.f2h_RREADY         (),                                //                  .rready
		.h2f_lw_axi_clk     (sys_sdram_pll_0_sys_clk_clk),     //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID        (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR      (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN       (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE      (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST     (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK      (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE     (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT      (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID     (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY     (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID         (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA       (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB       (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST       (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID      (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY      (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID         (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP       (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID      (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY      (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID        (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR      (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN       (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE      (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST     (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK      (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE     (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT      (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID     (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY     (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID         (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA       (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP       (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST       (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID      (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY      (hps_0_h2f_lw_axi_master_rready)   //                  .rready
	);

	DE1_SOC_jtag_uart_0 jtag_uart_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                                 //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         ()                                                             //               irq.irq
	);

	single_port_ram #(
		.DATA_WIDTH (8),
		.ADDR_WIDTH (6)
	) single_port_ram_0 (
		.data    (mm_interconnect_0_single_port_ram_0_avalon_slave_0_writedata), // avalon_slave_0.writedata
		.addr    (mm_interconnect_0_single_port_ram_0_avalon_slave_0_address),   //               .address
		.we      (mm_interconnect_0_single_port_ram_0_avalon_slave_0_write),     //               .write
		.q       (mm_interconnect_0_single_port_ram_0_avalon_slave_0_readdata),  //               .readdata
		.clk     (sys_sdram_pll_0_sys_clk_clk),                                  //          clock.clk
		.reset_n (~rst_controller_reset_out_reset)                               //          reset.reset_n
	);

	DE1_SOC_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (clk_clk),                       //      ref_clk.clk
		.ref_reset_reset    (~hps_0_h2f_reset_reset),        //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk),   //      sys_clk.clk
		.sdram_clk_clk      (sys_sdram_pll_0_sdram_clk_clk), //    sdram_clk.clk
		.reset_source_reset ()                               // reset_source.reset
	);

	DE1_SOC_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                           (hps_0_h2f_axi_master_awid),                                    //                          hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                         (hps_0_h2f_axi_master_awaddr),                                  //                                              .awaddr
		.hps_0_h2f_axi_master_awlen                          (hps_0_h2f_axi_master_awlen),                                   //                                              .awlen
		.hps_0_h2f_axi_master_awsize                         (hps_0_h2f_axi_master_awsize),                                  //                                              .awsize
		.hps_0_h2f_axi_master_awburst                        (hps_0_h2f_axi_master_awburst),                                 //                                              .awburst
		.hps_0_h2f_axi_master_awlock                         (hps_0_h2f_axi_master_awlock),                                  //                                              .awlock
		.hps_0_h2f_axi_master_awcache                        (hps_0_h2f_axi_master_awcache),                                 //                                              .awcache
		.hps_0_h2f_axi_master_awprot                         (hps_0_h2f_axi_master_awprot),                                  //                                              .awprot
		.hps_0_h2f_axi_master_awvalid                        (hps_0_h2f_axi_master_awvalid),                                 //                                              .awvalid
		.hps_0_h2f_axi_master_awready                        (hps_0_h2f_axi_master_awready),                                 //                                              .awready
		.hps_0_h2f_axi_master_wid                            (hps_0_h2f_axi_master_wid),                                     //                                              .wid
		.hps_0_h2f_axi_master_wdata                          (hps_0_h2f_axi_master_wdata),                                   //                                              .wdata
		.hps_0_h2f_axi_master_wstrb                          (hps_0_h2f_axi_master_wstrb),                                   //                                              .wstrb
		.hps_0_h2f_axi_master_wlast                          (hps_0_h2f_axi_master_wlast),                                   //                                              .wlast
		.hps_0_h2f_axi_master_wvalid                         (hps_0_h2f_axi_master_wvalid),                                  //                                              .wvalid
		.hps_0_h2f_axi_master_wready                         (hps_0_h2f_axi_master_wready),                                  //                                              .wready
		.hps_0_h2f_axi_master_bid                            (hps_0_h2f_axi_master_bid),                                     //                                              .bid
		.hps_0_h2f_axi_master_bresp                          (hps_0_h2f_axi_master_bresp),                                   //                                              .bresp
		.hps_0_h2f_axi_master_bvalid                         (hps_0_h2f_axi_master_bvalid),                                  //                                              .bvalid
		.hps_0_h2f_axi_master_bready                         (hps_0_h2f_axi_master_bready),                                  //                                              .bready
		.hps_0_h2f_axi_master_arid                           (hps_0_h2f_axi_master_arid),                                    //                                              .arid
		.hps_0_h2f_axi_master_araddr                         (hps_0_h2f_axi_master_araddr),                                  //                                              .araddr
		.hps_0_h2f_axi_master_arlen                          (hps_0_h2f_axi_master_arlen),                                   //                                              .arlen
		.hps_0_h2f_axi_master_arsize                         (hps_0_h2f_axi_master_arsize),                                  //                                              .arsize
		.hps_0_h2f_axi_master_arburst                        (hps_0_h2f_axi_master_arburst),                                 //                                              .arburst
		.hps_0_h2f_axi_master_arlock                         (hps_0_h2f_axi_master_arlock),                                  //                                              .arlock
		.hps_0_h2f_axi_master_arcache                        (hps_0_h2f_axi_master_arcache),                                 //                                              .arcache
		.hps_0_h2f_axi_master_arprot                         (hps_0_h2f_axi_master_arprot),                                  //                                              .arprot
		.hps_0_h2f_axi_master_arvalid                        (hps_0_h2f_axi_master_arvalid),                                 //                                              .arvalid
		.hps_0_h2f_axi_master_arready                        (hps_0_h2f_axi_master_arready),                                 //                                              .arready
		.hps_0_h2f_axi_master_rid                            (hps_0_h2f_axi_master_rid),                                     //                                              .rid
		.hps_0_h2f_axi_master_rdata                          (hps_0_h2f_axi_master_rdata),                                   //                                              .rdata
		.hps_0_h2f_axi_master_rresp                          (hps_0_h2f_axi_master_rresp),                                   //                                              .rresp
		.hps_0_h2f_axi_master_rlast                          (hps_0_h2f_axi_master_rlast),                                   //                                              .rlast
		.hps_0_h2f_axi_master_rvalid                         (hps_0_h2f_axi_master_rvalid),                                  //                                              .rvalid
		.hps_0_h2f_axi_master_rready                         (hps_0_h2f_axi_master_rready),                                  //                                              .rready
		.sys_sdram_pll_0_sys_clk_clk                         (sys_sdram_pll_0_sys_clk_clk),                                  //                       sys_sdram_pll_0_sys_clk.clk
		.single_port_ram_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // single_port_ram_0_reset_reset_bridge_in_reset.reset
		.single_port_ram_0_avalon_slave_0_address            (mm_interconnect_0_single_port_ram_0_avalon_slave_0_address),   //              single_port_ram_0_avalon_slave_0.address
		.single_port_ram_0_avalon_slave_0_write              (mm_interconnect_0_single_port_ram_0_avalon_slave_0_write),     //                                              .write
		.single_port_ram_0_avalon_slave_0_readdata           (mm_interconnect_0_single_port_ram_0_avalon_slave_0_readdata),  //                                              .readdata
		.single_port_ram_0_avalon_slave_0_writedata          (mm_interconnect_0_single_port_ram_0_avalon_slave_0_writedata)  //                                              .writedata
	);

	DE1_SOC_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                  (hps_0_h2f_lw_axi_master_awid),                                //                 hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                (hps_0_h2f_lw_axi_master_awaddr),                              //                                        .awaddr
		.hps_0_h2f_lw_axi_master_awlen                 (hps_0_h2f_lw_axi_master_awlen),                               //                                        .awlen
		.hps_0_h2f_lw_axi_master_awsize                (hps_0_h2f_lw_axi_master_awsize),                              //                                        .awsize
		.hps_0_h2f_lw_axi_master_awburst               (hps_0_h2f_lw_axi_master_awburst),                             //                                        .awburst
		.hps_0_h2f_lw_axi_master_awlock                (hps_0_h2f_lw_axi_master_awlock),                              //                                        .awlock
		.hps_0_h2f_lw_axi_master_awcache               (hps_0_h2f_lw_axi_master_awcache),                             //                                        .awcache
		.hps_0_h2f_lw_axi_master_awprot                (hps_0_h2f_lw_axi_master_awprot),                              //                                        .awprot
		.hps_0_h2f_lw_axi_master_awvalid               (hps_0_h2f_lw_axi_master_awvalid),                             //                                        .awvalid
		.hps_0_h2f_lw_axi_master_awready               (hps_0_h2f_lw_axi_master_awready),                             //                                        .awready
		.hps_0_h2f_lw_axi_master_wid                   (hps_0_h2f_lw_axi_master_wid),                                 //                                        .wid
		.hps_0_h2f_lw_axi_master_wdata                 (hps_0_h2f_lw_axi_master_wdata),                               //                                        .wdata
		.hps_0_h2f_lw_axi_master_wstrb                 (hps_0_h2f_lw_axi_master_wstrb),                               //                                        .wstrb
		.hps_0_h2f_lw_axi_master_wlast                 (hps_0_h2f_lw_axi_master_wlast),                               //                                        .wlast
		.hps_0_h2f_lw_axi_master_wvalid                (hps_0_h2f_lw_axi_master_wvalid),                              //                                        .wvalid
		.hps_0_h2f_lw_axi_master_wready                (hps_0_h2f_lw_axi_master_wready),                              //                                        .wready
		.hps_0_h2f_lw_axi_master_bid                   (hps_0_h2f_lw_axi_master_bid),                                 //                                        .bid
		.hps_0_h2f_lw_axi_master_bresp                 (hps_0_h2f_lw_axi_master_bresp),                               //                                        .bresp
		.hps_0_h2f_lw_axi_master_bvalid                (hps_0_h2f_lw_axi_master_bvalid),                              //                                        .bvalid
		.hps_0_h2f_lw_axi_master_bready                (hps_0_h2f_lw_axi_master_bready),                              //                                        .bready
		.hps_0_h2f_lw_axi_master_arid                  (hps_0_h2f_lw_axi_master_arid),                                //                                        .arid
		.hps_0_h2f_lw_axi_master_araddr                (hps_0_h2f_lw_axi_master_araddr),                              //                                        .araddr
		.hps_0_h2f_lw_axi_master_arlen                 (hps_0_h2f_lw_axi_master_arlen),                               //                                        .arlen
		.hps_0_h2f_lw_axi_master_arsize                (hps_0_h2f_lw_axi_master_arsize),                              //                                        .arsize
		.hps_0_h2f_lw_axi_master_arburst               (hps_0_h2f_lw_axi_master_arburst),                             //                                        .arburst
		.hps_0_h2f_lw_axi_master_arlock                (hps_0_h2f_lw_axi_master_arlock),                              //                                        .arlock
		.hps_0_h2f_lw_axi_master_arcache               (hps_0_h2f_lw_axi_master_arcache),                             //                                        .arcache
		.hps_0_h2f_lw_axi_master_arprot                (hps_0_h2f_lw_axi_master_arprot),                              //                                        .arprot
		.hps_0_h2f_lw_axi_master_arvalid               (hps_0_h2f_lw_axi_master_arvalid),                             //                                        .arvalid
		.hps_0_h2f_lw_axi_master_arready               (hps_0_h2f_lw_axi_master_arready),                             //                                        .arready
		.hps_0_h2f_lw_axi_master_rid                   (hps_0_h2f_lw_axi_master_rid),                                 //                                        .rid
		.hps_0_h2f_lw_axi_master_rdata                 (hps_0_h2f_lw_axi_master_rdata),                               //                                        .rdata
		.hps_0_h2f_lw_axi_master_rresp                 (hps_0_h2f_lw_axi_master_rresp),                               //                                        .rresp
		.hps_0_h2f_lw_axi_master_rlast                 (hps_0_h2f_lw_axi_master_rlast),                               //                                        .rlast
		.hps_0_h2f_lw_axi_master_rvalid                (hps_0_h2f_lw_axi_master_rvalid),                              //                                        .rvalid
		.hps_0_h2f_lw_axi_master_rready                (hps_0_h2f_lw_axi_master_rready),                              //                                        .rready
		.sys_sdram_pll_0_sys_clk_clk                   (sys_sdram_pll_0_sys_clk_clk),                                 //                 sys_sdram_pll_0_sys_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // jtag_uart_0_reset_reset_bridge_in_reset.reset
		.jtag_uart_0_avalon_jtag_slave_address         (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //           jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write           (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_0_avalon_jtag_slave_read            (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_0_avalon_jtag_slave_readdata        (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata       (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect      (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect)   //                                        .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
