module matrix_ingest 
#(parameter DATA_WIDTH=64, parameter ADDR_WIDTH=1)
(
	input [(DATA_WIDTH-1):0] data,
	input [(ADDR_WIDTH-1):0] addr,
	input we, clk, reset_n,
	output [(DATA_WIDTH-1):0] q
);
	

	reg [DATA_WIDTH-1:0] ram[2**ADDR_WIDTH-1:0];

	// Variable to hold the registered read address
	reg [ADDR_WIDTH-1:0] addr_reg;
	
	mul_add_96 u0 (
		.data_in (data),
		.z (q)
	);
	
	
	always @ (posedge clk or negedge reset_n)
	begin
		if (!reset_n) begin
			addr_reg <= {ADDR_WIDTH{1'b0}};
		end
		// Write
		else begin
			if (we) begin
				ram[addr] <= data;
			addr_reg <= addr;
			end
		end
	end

endmodule 