module adb_populater (

);

endmodule
