module requester_weights
#(parameter num_engines=10)
(		
		//axi variables
		input [(DATA_WIDTH-1):0] data,
		input [(ADDR_WIDTH-1):0] addr,
		input we, clk, reset_n,
		output [(DATA_WIDTH-1):0] q,
		
		//info from and to engines:
		input  wire [num_engines-1:0] data_in,
		output wire [33:0] request
);




endmodule
